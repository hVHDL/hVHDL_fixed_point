-- intentionally empty, remove!

