library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;

package multiplier_pipeline_registers_pkg is

    constant input_registers  : integer := 1;
    constant output_registers : integer := 1;

end package multiplier_pipeline_registers_pkg;
